// https://github.com/balanx/LogicDesignLib

`ifndef  LDL_RTL_DEFINE_VH
`define  LDL_RTL_DEFINE_VH

`define  LDL_ALWAYS_STATEMENT(CLOCK, RESET)    \
    always @(posedge CLOCK, posedge RESET)

`endif // LDL_RTL_DEFINE_VH

// LDL.

