// https://github.com/balanx/LogicDesignLib

`ifndef  LDL_MACROS_VH
`define  LDL_MACROS_VH

`define  LDL_ALWAYS     \
    always @(posedge clk)

`endif // LDL_MACROS_VH

// LDL.

