// https://github.com/balanx/LogicDesignLib

`ifndef  LDL_MACROS_VH
`define  LDL_MACROS_VH

`define  LDL_ALWAYS_STATEMENT(CLOCK, RESET)    \
    always @(posedge CLOCK, posedge RESET)

`endif // LDL_MACROS_VH

// LDL.

